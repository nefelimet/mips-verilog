`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   18:52:01 01/17/2022
// Design Name:   PROCESSOR
// Module Name:   C:/Users/Nefel/Desktop/University/project1/PROCESSOR_tb.v
// Project Name:  project1
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: PROCESSOR
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module PROCESSOR_tb;

	// Inputs
	reg clk = 0;

	// Outputs
	wire [31:0] Instr;
	wire [31:0] Immed;
	wire [31:0] RF_A;
	wire [31:0] RF_B_or_sb;
	wire [31:0] ALU_out;
	wire [31:0] MEM_out;
	wire [31:0] lui_out;
	  
	// Instantiate the Unit Under Test (UUT)
	PROCESSOR uut (
		.clk(clk),
		.Instr(Instr),
		.Immed(Immed),
		.RF_A(RF_A),
		.RF_B_or_sb(RF_B_or_sb),
		.ALU_out(ALU_out),
		.MEM_out(MEM_out),
		.lui_out(lui_out)
	);

	always #1 clk = ~clk;

	initial begin
		
		$display("PC_out: %b", uut.if_stage.progcount.Dout);
		#2;
		$display("--------------1--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("PC_out: %b", uut.if_stage.progcount.Dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------2--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("PC_out: %b", uut.if_stage.progcount.Dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------3--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("PC_out: %b", uut.if_stage.progcount.Dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------4--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("PC_out: %b", uut.if_stage.progcount.Dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------5--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("PC_out: %b", uut.if_stage.progcount.Dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------6--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------7--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------8--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------9--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------10--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------11--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------12--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------13--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------14--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------15--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------16--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------17--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------18--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("PC_out: %b", uut.if_stage.progcount.Dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------19--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("PC_out: %b", uut.if_stage.progcount.Dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------20--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("PC_out: %b", uut.if_stage.progcount.Dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------21--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("PC_out: %b", uut.if_stage.progcount.Dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------22--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("PC_out: %b", uut.if_stage.progcount.Dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------23--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("PC_out: %b", uut.if_stage.progcount.Dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------24--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("PC_out: %b", uut.if_stage.progcount.Dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------25--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("PC_out: %b", uut.if_stage.progcount.Dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------26--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("PC_out: %b", uut.if_stage.progcount.Dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------27--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("PC_out: %b", uut.if_stage.progcount.Dout);
		$display("-----------------------------");
		
		#2;
		//sw
		$display("--------------28--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("MEM addr: %b, MEM Din: %b, MEM WrEn: %b, MEM Dout: %b", uut.mem_stage.ram_mem.addr, uut.mem_stage.ram_mem.din, uut.mem_stage.ram_mem.we, uut.mem_stage.ram_mem.dout);
		$display("RF_B: %b, sb_out: %b, RF_B_or_sb: %b", uut.dec_stage.RF.r5.Dout, uut.dec_stage.sb_out, uut.dec_stage.RF_B_or_sb);
		$display("PC_out: %b", uut.if_stage.progcount.Dout);
		$display("-----------------------------");
		
		#2;
		//sb
		$display("--------------29--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("MEM addr: %b, MEM Din: %b, MEM WrEn: %b, MEM Dout: %b", uut.mem_stage.ram_mem.addr, uut.mem_stage.ram_mem.din, uut.mem_stage.ram_mem.we, uut.mem_stage.ram_mem.dout);
		$display("RF_B: %b, sb_out: %b, RF_B_or_sb: %b", uut.dec_stage.RF.r10.Dout, uut.dec_stage.sb_out, uut.dec_stage.RF_B_or_sb);
		$display("-----------------------------");
		
		#2;
		$display("--------------30--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("MEM addr: %b, MEM Din: %b, MEM WrEn: %b, MEM Dout: %b", uut.mem_stage.ram_mem.addr, uut.mem_stage.ram_mem.din, uut.mem_stage.ram_mem.we, uut.mem_stage.ram_mem.dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------31--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("MEM addr: %b, MEM Din: %b, MEM WrEn: %b, MEM Dout: %b", uut.mem_stage.ram_mem.addr, uut.mem_stage.ram_mem.din, uut.mem_stage.ram_mem.we, uut.mem_stage.ram_mem.dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------32--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("MEM addr: %b, MEM Din: %b, MEM WrEn: %b, MEM Dout: %b", uut.mem_stage.ram_mem.addr, uut.mem_stage.ram_mem.din, uut.mem_stage.ram_mem.we, uut.mem_stage.ram_mem.dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------33--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("MEM addr: %b, MEM Din: %b, MEM WrEn: %b, MEM Dout: %b", uut.mem_stage.ram_mem.addr, uut.mem_stage.ram_mem.din, uut.mem_stage.ram_mem.we, uut.mem_stage.ram_mem.dout);
		$display("-----------------------------");
		
		#2;
		$display("--------------34--------------");
		$display("Instr = %b", uut.Instr);
		$display("PC_sel = %b, PC_LdEn = %b, RF_WrEn = %b, RF_WrData_sel = %b, RF_B_sel = %b", uut.PC_sel, uut.PC_LdEn, uut.RF_WrEn, uut.RF_WrData_sel, uut.RF_B_sel);
		$display("ALU_Bin_sel = %b, ALU_func = %b, Mem_WrEn = %b, lui = %b, lb = %b, sb = %b", uut.ALU_Bin_sel, uut.ALU_func, uut.Mem_WrEn, uut.lui, uut.lb, uut.sb);
		$display("RF_A = %b, RF_B_or_sb = %b, Immed = %b, ALU_out = %b", uut.RF_A, uut.RF_B_or_sb, uut.Immed, uut.ALU_out);
		$display("r0 Dout: %b", uut.dec_stage.RF.r0.Dout);
		$display("r1 Dout: %b", uut.dec_stage.RF.r1.Dout);
		$display("r2 Dout: %b", uut.dec_stage.RF.r2.Dout);
		$display("r3 Dout: %b", uut.dec_stage.RF.r3.Dout);
		$display("r4 Dout: %b", uut.dec_stage.RF.r4.Dout);
		$display("r5 Dout: %b", uut.dec_stage.RF.r5.Dout);
		$display("r6 Dout: %b", uut.dec_stage.RF.r6.Dout);
		$display("r7 Dout: %b", uut.dec_stage.RF.r7.Dout);
		$display("r8 Dout: %b", uut.dec_stage.RF.r8.Dout);
		$display("r9 Dout: %b", uut.dec_stage.RF.r9.Dout);
		$display("r10 Dout: %b", uut.dec_stage.RF.r10.Dout);
		$display("r11 Dout: %b", uut.dec_stage.RF.r11.Dout);
		$display("r12 Dout: %b", uut.dec_stage.RF.r12.Dout);
		$display("r13 Dout: %b", uut.dec_stage.RF.r13.Dout);
		$display("r14 Dout: %b", uut.dec_stage.RF.r14.Dout);
		$display("r15 Dout: %b", uut.dec_stage.RF.r15.Dout);
		$display("r16 Dout: %b", uut.dec_stage.RF.r16.Dout);
		$display("r17 Dout: %b", uut.dec_stage.RF.r17.Dout);
		$display("r18 Dout: %b", uut.dec_stage.RF.r18.Dout);
		$display("r19 Dout: %b", uut.dec_stage.RF.r19.Dout);
		$display("r20 Dout: %b", uut.dec_stage.RF.r20.Dout);
		$display("r21 Dout: %b", uut.dec_stage.RF.r21.Dout);
		$display("r22 Dout: %b", uut.dec_stage.RF.r22.Dout);
		$display("r23 Dout: %b", uut.dec_stage.RF.r23.Dout);
		$display("r24 Dout: %b", uut.dec_stage.RF.r24.Dout);
		$display("r25 Dout: %b", uut.dec_stage.RF.r25.Dout);
		$display("r26 Dout: %b", uut.dec_stage.RF.r26.Dout);
		$display("r27 Dout: %b", uut.dec_stage.RF.r27.Dout);
		$display("r28 Dout: %b", uut.dec_stage.RF.r28.Dout);
		$display("r29 Dout: %b", uut.dec_stage.RF.r29.Dout);
		$display("r30 Dout: %b", uut.dec_stage.RF.r30.Dout);
		$display("r31 Dout: %b", uut.dec_stage.RF.r31.Dout);
		$display("instr2: %b, read_reg2: %b, RF_B: %b", uut.dec_stage.instr2, uut.dec_stage.read_reg2, uut.dec_stage.RF.Dout2);
		$display("MEM: %b", uut.mem_stage.ram_mem.dout);
		$display("MEM addr: %b, MEM Din: %b, MEM WrEn: %b, MEM Dout: %b", uut.mem_stage.ram_mem.addr, uut.mem_stage.ram_mem.din, uut.mem_stage.ram_mem.we, uut.mem_stage.ram_mem.dout);
		$display("-----------------------------");
		
	//Simulation time: 34*2=68ns
	end
      
endmodule

